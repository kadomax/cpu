
//opcodes
`define ADD_OPCODE 4'b0000
`define SUB_OPCODE 4'b0001
`define AND_OPCODE 4'b0010
`define OR_OPCODE 4'b0011
`define XOR_OPCODE 4'b0010
`define B_OPCODE 4'b0101
`define BP_OPCODE 4'b0110
`define BN_OPCODE 4'b0111
`define BZ_OPCODE 4'b1000
`define LDRIA_OPCODE 4'b1001
`define LDRIB_OPCODE 4'b1010
`define LDRA_OPCODE 4'b1011
`define LDRB_OPCODE 4'b1100
`define STR_OPCODE 4'b1101
`define NOP_OPCODE 4'b1110
`define HLT_OPCODE 4'b1111